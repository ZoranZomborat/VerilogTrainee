library verilog;
use verilog.vl_types.all;
entity func is
end func;
